library ieee ;
	use ieee.std_logic_1164.all ;
	use ieee.numeric_std.all ;

entity TDESStateMachine is
  port (
	clock : IN STD_LOGIC;
	done : OUT STD_LOGIC;
  ) ;
end entity ; -- TDESStateMachine

architecture arch of TDESStateMachine is

begin

end architecture ; -- arch