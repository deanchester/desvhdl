library ieee ;
	use ieee.std_logic_1164.all ;
	use ieee.numeric_std.all ;

entity CryptoCore is
  port (
	clock
  ) ;
end entity ; -- CryptoCore

architecture arch of CryptoCore is

begin

end architecture ; -- arch